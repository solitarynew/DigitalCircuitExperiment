module block();


endmodule
