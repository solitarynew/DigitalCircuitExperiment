module decode_hex(count,);