module unblock();


endmodule
